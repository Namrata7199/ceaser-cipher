module Verilog_BM_121_202(input a,input b,input c,input d,input e,input f,input g,input h,input i,input j,input k,input l,input m,input n,input o,input p,input q,input r,input s,input t,input u,input v,input w,input x,input y,input z,input i1,input i2,input i3,input i4,input i5,input i6,input i7,input i8,input i9,input i10,input i11,input i12,input i13,input i14,input i15,input i16,input i17,input i18,input i19,input i20,input i21,input i22,input i23,input i24,input i25,input i26,input en,input cap,output reg [7:0]out);
reg [4:0]w1;
reg [4:0]w2;
reg [5:0]w3;
reg [5:0]s0;
reg [5:0]w4;
reg [6:0]w5;
reg [6:0]s1;
reg [6:0]w6;
reg [7:0]s2;
integer x0;
always@(*)
begin
	if(a==1)
		w1=0;
	if(b==1)
		w1=1;
	if(c==1)
		w1=2;
	if(d==1)
		w1=3;
	if(e==1)
		w1=4;
	if(f==1)
		w1=5;
	if(g==1)
		w1=6;
	if(h==1)
		w1=7;
	if(i==1)
		w1=8;
	if(j==1)
		w1=9;
	if(k==1)
		w1=10;
	if(l==1)
		w1=11;
	if(m==1)
		w1=12;
	if(n==1)
		w1=13;
	if(o==1)
		w1=14;
	if(p==1)
		w1=15;
	if(q==1)
		w1=16;
	if(r==1)
		w1=17;
	if(s==1)
		w1=18;
	if(t==1)
		w1=19;
	if(u==1)
		w1=20;
	if(v==1)
		w1=21;
	if(w==1)
		w1=22;
	if(x==1)
		w1=23;
	if(y==1)
		w1=24;
	if(z==1)
		w1=25;
	if(i1==1)
		w2=1;
	if(i2==1)
		w2=2;
	if(i3==1)
		w2=3;
	if(i4==1)
		w2=4;
	if(i5==1)
		w2=5;
	if(i6==1)
		w2=6;
	if(i7==1)
		w2=7;
	if(i8==1)
		w2=8;
	if(i9==1)
		w2=9;
	if(i10==1)
		w2=10;
	if(i11==1)
		w2=11;
	if(i12==1)
		w2=12;
	if(i13==1)
		w2=13;
	if(i14==1)
		w2=14;
	if(i15==1)
		w2=15;
	if(i16==1)
		w2=16;
	if(i17==1)
		w2=17;
	if(i18==1)
		w2=18;
	if(i19==1)
		w2=19;
	if(i20==1)
		w2=20;
	if(i21==1)
		w2=21;
	if(i22==1)
		w2=22;
	if(i23==1)
		w2=23;
	if(i24==1)
		w2=24;
	if(i25==1)
		w2=25;
	if(i26==1)
		w2=26;
	for(x0=0;x0<5;x0=x0+1)
	begin
		w2[x0]=w2[x0]^en;
	end
	s0[0]=en;
	for(x0=0;x0<5;x0=x0+1)
	begin
		w3[x0]=s0[x0]^w1[x0]^w2[x0];
		s0[x0+1]=(s0[x0]&w1[x0])|(s0[x0]&w2[x0])|(w1[x0]&w2[x0]);
	end
	w3[5]=s0[5];
	if(w3>=6'b011010||w3<6'b000000)
	begin
		if(en==0)
		begin
			w4=6'b100101;
		end
		else
		begin
			w4=6'b011010;
		end
		s1[0]=~en;
		for(x0=0;x0<6;x0=x0+1)
		begin
			w5[x0]=s1[x0]^w3[x0]^w4[x0];
			s1[x0+1]=(s1[x0]&w3[x0])|(s1[x0]&w4[x0])|(w3[x0]&w4[x0]);
		end
		w5[6]=s1[6];
	end
	else
	begin
		for(x0=0;x0<6;x0=x0+1)
		begin
			w5[x0]=w3[x0];
		end
		w5[6]=0;
	end
	if(cap==0)
		w6=97;
	else w6=65;
	s2[0]=1'b0;
	for(x0=0;x0<7;x0=x0+1)
	begin
		out[x0]=s2[x0]^w6[x0]^w5[x0];
		s2[x0+1]=(s2[x0]&w6[x0])|(s2[x0]&w5[x0])|(w5[x0]&w6[x0]);
	end
	out[7]=s2[7];
end
endmodule
